module display(sec, min, hour, day, mont, year,a,b,c,d,e,f,g);
    input [5:0]	sec;
	input [5:0]	min;
	input [4:0]	hour;
	input [4:0]	day;
	input [3:0]	mont;
	input [12:0] year;
    output [13:0] a,b,c,d,e,f,g;
    
    wire [3:0] sec_0,sec_1,min_0,min_1,hour_0,hour_1,day_0,day_1,mont_0,mont_1,year_0,year_1,year_2,year_3;
    assign sec_0=sec%10;
    assign sec_1=sec/10;
    assign min_0=min%10;
    assign min_1=min/10;
    assign hour_0=hour%10;
    assign hour_1=hour/10;
    assign day_0=day%10;
    assign day_1=day/10;
    assign mont_0=mont%10;
    assign mont_1=mont/10;
    assign year_0=year%10;
    assign year_1=((year-year_0)/10)%10;
    assign year_2=((year-year_0-year_1*10)/100)%10;
    assign year_3=year/1000;
    
    giaima7thanh m_0    (.x(sec_0),.a(a[0]),.b(b[0]),.c(c[0]),.d(d[0]),.e(e[0]),.f(f[0]),.g(g[0]));
    giaima7thanh m_1    (.x(sec_1),.a(a[1]),.b(b[1]),.c(c[1]),.d(d[1]),.e(e[1]),.f(f[1]),.g(g[1]));
    giaima7thanh m_2    (.x(min_0),.a(a[2]),.b(b[2]),.c(c[2]),.d(d[2]),.e(e[2]),.f(f[2]),.g(g[2]));
    giaima7thanh m_3    (.x(min_1),.a(a[3]),.b(b[3]),.c(c[3]),.d(d[3]),.e(e[3]),.f(f[3]),.g(g[3]));
    giaima7thanh m_4    (.x(hour_0),.a(a[4]),.b(b[4]),.c(c[4]),.d(d[4]),.e(e[4]),.f(f[4]),.g(g[4]));
    giaima7thanh m_5    (.x(hour_1),.a(a[5]),.b(b[5]),.c(c[5]),.d(d[5]),.e(e[5]),.f(f[5]),.g(g[5]));
    giaima7thanh m_6    (.x(day_0),.a(a[6]),.b(b[6]),.c(c[6]),.d(d[6]),.e(e[6]),.f(f[6]),.g(g[6]));
    giaima7thanh m_7    (.x(day_1),.a(a[7]),.b(b[7]),.c(c[7]),.d(d[7]),.e(e[7]),.f(f[7]),.g(g[7]));
    giaima7thanh m_8    (.x(mont_0),.a(a[8]),.b(b[8]),.c(c[8]),.d(d[8]),.e(e[8]),.f(f[8]),.g(g[8]));
    giaima7thanh m_9    (.x(mont_1),.a(a[9]),.b(b[9]),.c(c[9]),.d(d[9]),.e(e[9]),.f(f[9]),.g(g[9]));
    giaima7thanh m_10   (.x(year_0),.a(a[10]),.b(b[10]),.c(c[10]),.d(d[10]),.e(e[10]),.f(f[10]),.g(g[10]));
    giaima7thanh m_11   (.x(year_1),.a(a[11]),.b(b[11]),.c(c[11]),.d(d[11]),.e(e[11]),.f(f[11]),.g(g[11]));
    giaima7thanh m_12   (.x(year_2),.a(a[12]),.b(b[12]),.c(c[12]),.d(d[12]),.e(e[12]),.f(f[12]),.g(g[12]));
    giaima7thanh m_13   (.x(year_3),.a(a[13]),.b(b[13]),.c(c[13]),.d(d[13]),.e(e[13]),.f(f[13]),.g(g[13]));
endmodule
